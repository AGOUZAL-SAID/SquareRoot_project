library ieee ;
use ieee.std_logic_1164.all ;
use ieee.numeric_std.all ;



entity TB_AV is
    generic(NBITS : integer := 32) ;
end entity;

architecture a1 of TB_AV is
begin 
end a1;