library ieee ;
use ieee.std_logic_1164.all ;
use ieee.numeric_std.all ;



entity TB_INST is
end entity;

architecture a1 of TB_INST is
begin 
-- Nothing for the moment 
end a1;